gp_pos_cam_inst : gp_pos_cam PORT MAP (
		pattern	 => pattern_sig,
		wraddress	 => wraddress_sig,
		wren	 => wren_sig,
		inclock	 => inclock_sig,
		mbits	 => mbits_sig
	);
