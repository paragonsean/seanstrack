------------------- QUAD_DECODER.VHD ------------------------
----------- Copyright 2002, Visi-Trak Worldwide -------------
--
-- 2-8-02 This version of quad decoder outputs 4 speed pulses, 1 for each
-- of the quadrature quadrants.  If interfacing to a standard single 
-- quadrant velocity circuit, use the speed_pulse_main output as the speed pulse.


-- 10-2-02 Elminated speed_pulse_main.  Speed pulses are now simply
-- speed_pulse_q1,2,3 and 4. 
-- When moving forward, the quadrants are defined as follows:
-- 		Q1 --> Rise to rise, chA
--		Q2 --> Rise to rise, chB
--		Q3 --> Fall to fall, chA
--		Q4 --> Fall to fall, chB
-- When moving in reverse, the quadrants are defined as follows:
-- 		Q4 --> Rise to rise, chB
--		Q3 --> Rise to rise, chA
--		Q2 --> Fall to fall, chB
--		Q1 --> Fall to fall, chA
-- The speed pulses are now directly generated by the edges as just 
-- defined.  Perviously they were generated by a counter keeping track
-- of X4 pulses.  There was no way to definitively link a given speed 
-- pulse with a specific quadrant.  Now there is.
--
-- When a quadrature error or up/down change is detected, once direction
-- change is established, the next 4 X4 counts will not generate speed
-- pulses.  After this, the next 4 speed pulses generated will have either
-- the UD changed or quad error bit set to allow marking the latched data
-- accordingly.  This will flag that data so the software can take the 
-- appropriate steps.


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


entity quad_decoder is
	port(
		clk			: in	std_logic;
		rst			: in	std_logic;  
		ch_a		: in	std_logic;
		ch_b		: in	std_logic;
		ch_a_out	: out	std_logic;	 	-- Registered ch_a
		ch_b_out	: out	std_logic;  	-- Registered ch_b
		speed_pulse_q1	: out	std_logic;	-- Must update speed pulse if up_dn changes a'la Prince
		speed_pulse_q2	: out	std_logic;
		speed_pulse_q3	: out	std_logic;
		speed_pulse_q4 : out	std_logic; 
		up_dn		: out 	std_logic;
		x4			: out	std_logic;
		up_dn_changed_out : out std_logic;
		err			: out	std_logic); 
end quad_decoder;


architecture behave OF quad_decoder is

signal CNT : std_logic_vector(2 downto 0);
signal UP_DN_CHANGED, LATCHED_UP_DN_CHANGED : std_logic;
signal RAW_SP_Q1, RAW_SP_Q2, RAW_SP_Q3, RAW_SP_Q4 : std_logic;
signal X4_INTERNAL, UP_DN_INTERNAL : std_logic;
signal AAA, BBB, TMPAA, TMPBB : std_logic;
signal QUADRATURE_ERROR, LATCHED_QUADRATURE_ERROR : std_logic;
signal REQUEST_FOR_SP_Q1, REQUEST_FOR_SP_Q2 : std_logic;
signal REQUEST_FOR_SP_Q3, REQUEST_FOR_SP_Q4 : std_logic;
signal OK_TO_REMOVE_UD_CHANGED, OK_TO_REMOVE_QUADRATURE_ERROR : std_logic;

begin
-- This version of quadrature decoder is completely syncronous in operation.



-- This process keeps track of x4 counts after a reset or after a change
-- in up/down or after a quadrature error.  Speed pulses will be inhibited
-- until four X4 counts have occured after one of the above conditions.
-- CNT will count up to and stay at "101" until U/D changes or reset.
-- Once CNT reaches "101", five X4 counts will have beed counted.  
-- Speed pulses will be enabled on the 5th. X4 count received.
process (clk, rst)
		begin
		if rst = '1' or UP_DN_CHANGED = '1' or QUADRATURE_ERROR = '1' then
			CNT <= "000";
			
		elsif (clk 'event and clk = '1') then	
			if (X4_INTERNAL = '1' and UP_DN_INTERNAL = '1') then -- Remove UP_DN_INTERNAL condition to collect data in reverse
				
				-- CNT Stays at "111" until U/D changes, quad error or reset.
				if (CNT < "111") then				
				  CNT <= CNT + '1'; -- Only increment if moving forward.
				else null;
				end if;
					
			else null;
			end if;
		else null;
		end if;	
end process;




-- Process to process the UP_DN_CHANGED signal.  No need put rst in the
-- sensitivity list.  The quad decoder process will assert UP_DN_CHANGED
-- at reset.
process(clk)
	begin
	if (clk 'event and clk = '1') then
		OK_TO_REMOVE_UD_CHANGED <= '0';
		
		if (UP_DN_CHANGED = '1') then
			LATCHED_UP_DN_CHANGED <= '1';
		-- When the 8th. X4 pulse is counted, remove the U/D changed signal	
		elsif ((LATCHED_UP_DN_CHANGED = '1' and CNT = "111") and X4_INTERNAL = '1') then
			OK_TO_REMOVE_UD_CHANGED <= '1';
		elsif (OK_TO_REMOVE_UD_CHANGED = '1') then 
			LATCHED_UP_DN_CHANGED <= '0';
		else null;	
		end if;	
	else null;
	end if;
end process;

up_dn_changed_out <= LATCHED_UP_DN_CHANGED;


-- Process to process the QUADRATURE_ERROR signal.  
process(clk, rst)
	begin
	if (rst = '1') then
		LATCHED_QUADRATURE_ERROR <= '0';
		OK_TO_REMOVE_QUADRATURE_ERROR <= '0';
	elsif (clk 'event and clk = '1') then
		OK_TO_REMOVE_QUADRATURE_ERROR <= '0';
		
		if (QUADRATURE_ERROR = '1') then
			LATCHED_QUADRATURE_ERROR <= '1';
		-- When the 8th. X4 pulse is counted, remove the quad error signal	
		elsif ((LATCHED_QUADRATURE_ERROR = '1' and CNT = "111") and X4_INTERNAL = '1') then
			OK_TO_REMOVE_QUADRATURE_ERROR <= '1';
		elsif (OK_TO_REMOVE_QUADRATURE_ERROR = '1') then
			LATCHED_QUADRATURE_ERROR <= '0';
		else null;
		end if;	
	else null;
	end if;
end process;

err <= LATCHED_QUADRATURE_ERROR;



-- Quadrature decoder
--
-- The quadrature decoder will decode the channel A and B transducer pulses
-- and generate the necessary signals for connecting the decoder to the
-- position and velocity counter circuits.
process (clk, rst)
	variable STATE	: std_logic_vector (3 downto 0);
	variable CLK_CTR : std_logic_vector (1 downto 0);
	variable REQUEST_FOR_X4_PULSE, OK_FOR_X4_PULSE, PREV_UP_DN : std_logic;
	begin
		if (rst = '1') then  -- Async reset
			PREV_UP_DN := UP_DN_INTERNAL;
			REQUEST_FOR_X4_PULSE := '0';
			OK_FOR_X4_PULSE := '0';
			X4_INTERNAL <= '0';
			UP_DN_CHANGED <= '1';
			UP_DN_INTERNAL <= '1';
			AAA <= '0';
			BBB <= '0';
			TMPAA <= '0';
			TMPBB <= '0';
			STATE := "0000";
			REQUEST_FOR_SP_Q1 <= '0';
			REQUEST_FOR_SP_Q2 <= '0';
			REQUEST_FOR_SP_Q3 <= '0';
			REQUEST_FOR_SP_Q4 <= '0';
			QUADRATURE_ERROR <= '0';
			CLK_CTR := "00";
		elsif (clk 'event and clk = '1') then
		 	   AAA <= TMPAA; BBB <= TMPBB;		-- Preserve the current states
			   TMPAA <= ch_a; TMPBB <= ch_b;	-- And get the new states
			   STATE := BBB & AAA & TMPBB & TMPAA;	-- aaa and bbb previous ch_a and ch_b states, aa and bb are the current states
				
				X4_INTERNAL <= '0';	
				QUADRATURE_ERROR <= '0';
				
				-- Now process 4x pulse requests.  If up_dn has changed, hold
				-- another clock cycle to allow up_dn to settle.
				if (PREV_UP_DN /= UP_DN_INTERNAL) then
					UP_DN_CHANGED <= '1'; 
					PREV_UP_DN := UP_DN_INTERNAL;
				elsif (REQUEST_FOR_X4_PULSE = '1') then
					OK_FOR_X4_PULSE := '1';
					REQUEST_FOR_X4_PULSE := '0';
				elsif (OK_FOR_X4_PULSE = '1') then 	
					X4_INTERNAL <= '1';
					OK_FOR_X4_PULSE := '0';
					UP_DN_CHANGED <= '0';
				else null;
				end if;
				
				case STATE is
					-- CLK_CTR is reset every X4 count.  It is incremented
					-- every clk cycle.  By the time it gets to "11" it's
					-- safe to process another count state.  If another
					-- count state occurs before this counter reaches "11"
					-- this will be defined as a quadrature error.  The 
					-- edges are too close together.
					when "0001"=> -- Count up quadrant #1
						if (CLK_CTR < "11") then -- Recently processed an X4 count, must be a quad error!
							OK_FOR_X4_PULSE := '0';
							QUADRATURE_ERROR <= '1';
						else	
						    UP_DN_INTERNAL <= '1'; -- Active high for count up
							REQUEST_FOR_X4_PULSE := '1';
							REQUEST_FOR_SP_Q1 <= '1';
			            	REQUEST_FOR_SP_Q2 <= '0';
			            	REQUEST_FOR_SP_Q3 <= '0';
			            	REQUEST_FOR_SP_Q4 <= '0';
							CLK_CTR := "00";
						end if;
			        when "0111"=> -- Count up quadrant #2
						if (CLK_CTR < "11") then -- Recently processed an X4 count, must be a quad error!
							OK_FOR_X4_PULSE := '0';
							QUADRATURE_ERROR <= '1';
						else
							UP_DN_INTERNAL <= '1'; -- Active high for count up
							REQUEST_FOR_X4_PULSE := '1';
							REQUEST_FOR_SP_Q1 <= '0';
			            	REQUEST_FOR_SP_Q2 <= '1';
			            	REQUEST_FOR_SP_Q3 <= '0';
			            	REQUEST_FOR_SP_Q4 <= '0';
							CLK_CTR := "00";
						end if;
			        when "1110"=> -- Count up quadrant #3
						if (CLK_CTR < "11") then -- Recently processed an X4 count, must be a quad error!
							OK_FOR_X4_PULSE := '0';
							QUADRATURE_ERROR <= '1';
						else
							UP_DN_INTERNAL <= '1'; -- Active high for count up
							REQUEST_FOR_X4_PULSE := '1';
							REQUEST_FOR_SP_Q1 <= '0';
			            	REQUEST_FOR_SP_Q2 <= '0';
			            	REQUEST_FOR_SP_Q3 <= '1';
			            	REQUEST_FOR_SP_Q4 <= '0';
							CLK_CTR := "00";
						end if;
			        when "1000"=> -- Count up quadrant #4
						if (CLK_CTR < "11") then -- Recently processed an X4 count, must be a quad error!
							OK_FOR_X4_PULSE := '0';
							QUADRATURE_ERROR <= '1';
						else
							UP_DN_INTERNAL <= '1'; -- Active high for count up
							REQUEST_FOR_X4_PULSE := '1';
							REQUEST_FOR_SP_Q1 <= '0';
			            	REQUEST_FOR_SP_Q2 <= '0';
			            	REQUEST_FOR_SP_Q3 <= '0';
			            	REQUEST_FOR_SP_Q4 <= '1';
							CLK_CTR := "00";
						end if;
			        when "0010"=> -- Count down quadrant #4
						if (CLK_CTR < "11") then -- Recently processed an X4 count, must be a quad error!
							OK_FOR_X4_PULSE := '0';
							QUADRATURE_ERROR <= '1';
						else
							UP_DN_INTERNAL <= '0';
							REQUEST_FOR_X4_PULSE := '1';
							REQUEST_FOR_SP_Q1 <= '0';
			            	REQUEST_FOR_SP_Q2 <= '0';
			            	REQUEST_FOR_SP_Q3 <= '0';
			            	REQUEST_FOR_SP_Q4 <= '1';
							CLK_CTR := "00";
						end if;
			        when "1011"=> -- Count down quadrant #3
						if (CLK_CTR < "11") then -- Recently processed an X4 count, must be a quad error!
							OK_FOR_X4_PULSE := '0';
							QUADRATURE_ERROR <= '1';
						else
							UP_DN_INTERNAL <= '0';
							REQUEST_FOR_X4_PULSE := '1';
							REQUEST_FOR_SP_Q1 <= '0';
			            	REQUEST_FOR_SP_Q2 <= '0';
			            	REQUEST_FOR_SP_Q3 <= '1';
			            	REQUEST_FOR_SP_Q4 <= '0';
							CLK_CTR := "00";
						end if;
			        when "1101"=> -- Count down quadrant #2
						if (CLK_CTR < "11") then -- Recently processed an X4 count, must be a quad error!
							OK_FOR_X4_PULSE := '0';
							QUADRATURE_ERROR <= '1';
						else
							UP_DN_INTERNAL <= '0';
							REQUEST_FOR_X4_PULSE := '1';
							REQUEST_FOR_SP_Q1 <= '0';
			            	REQUEST_FOR_SP_Q2 <= '1';
			           	 	REQUEST_FOR_SP_Q3 <= '0';
			            	REQUEST_FOR_SP_Q4 <= '0';
							CLK_CTR := "00";
						end if;
			        when "0100"=> -- Count down quadrant #1
						if (CLK_CTR < "11") then -- Recently processed an X4 count, must be a quad error!
							OK_FOR_X4_PULSE := '0';
							QUADRATURE_ERROR <= '1';
						else
							UP_DN_INTERNAL <= '0';
							REQUEST_FOR_X4_PULSE := '1';
							REQUEST_FOR_SP_Q1 <= '1';
			            	REQUEST_FOR_SP_Q2 <= '0';
			            	REQUEST_FOR_SP_Q3 <= '0';
			            	REQUEST_FOR_SP_Q4 <= '0';
							CLK_CTR := "00";
						end if;
			        when "0011"|"0110"|"1001"|"1100"=> -- Error states
						QUADRATURE_ERROR <= '1';
						X4_INTERNAL <= '0';
						REQUEST_FOR_X4_PULSE := '0';
						
					when others=>
						null;
				end case;
				
				if (REQUEST_FOR_X4_PULSE = '0') then
					if (CLK_CTR < "11") then
						CLK_CTR := CLK_CTR + '1';
					else null;
					end if;	
				else null;
				end if;
		else null;
		end if;
end process;

x4 <= X4_INTERNAL;
up_dn <= UP_DN_INTERNAL;
ch_a_out <= TMPAA;
ch_b_out <= TMPBB;


process(clk,rst)
begin
if (rst = '1') then
	speed_pulse_q1 <= '0';
	speed_pulse_q2 <= '0';
	speed_pulse_q3 <= '0';
	speed_pulse_q4 <= '0';
elsif (clk 'event and clk = '1') then
	speed_pulse_q1 <= '0';
	speed_pulse_q2 <= '0';
	speed_pulse_q3 <= '0';
	speed_pulse_q4 <= '0';
	if (CNT >= "101") then
		if (REQUEST_FOR_SP_Q1 = '1') then
			speed_pulse_q1 <= '1';
		else null;
		end if;
		
		if (REQUEST_FOR_SP_Q2 = '1') then
			speed_pulse_q2 <= '1';
		else null;
		end if;
		
		if (REQUEST_FOR_SP_Q3 = '1') then
			speed_pulse_q3 <= '1';
		else null;
		end if;
		
		if (REQUEST_FOR_SP_Q4 = '1') then
			speed_pulse_q4 <= '1';
		else null;
		end if;	
	else null;
	end if;
else null;
end if;
end process;

end behave;



